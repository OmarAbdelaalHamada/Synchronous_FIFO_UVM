package shared_pkg;
parameter FIFO_WIDTH = 16;
parameter FIFO_DEPTH = 8;
integer RD_EN_ON_DIST = 30;
integer WR_EN_ON_DIST = 70;
endpackage